module CPU (input logic clk, reset, 
	 output logic [31:0] PCF, 
	 input logic [31:0] InstrF, 
	 output logic MemWriteM, 
	 output logic [31:0] ALUOutM, WriteDataM,
	 input logic [31:0] ReadDataM);
//Cables


//Controller
//Hazard
endmodule